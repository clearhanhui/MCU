library verilog;
use verilog.vl_types.all;
entity MCU_vlg_vec_tst is
end MCU_vlg_vec_tst;
